<<<<<<< HEAD
module PCadder(result, oldPC);
	input [31:0] oldPC;
	output [31:0] result;
	assign result = oldPC + 4;
endmodule
=======
module PCadder(resultd, oldPC);
	input [31:0] oldPC;
	output [31:0] resultd;
	assign resultd = oldPC + 4;
endmodule
>>>>>>> 14f980056707609f192789c3457eade4c2ae4280
